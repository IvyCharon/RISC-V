`include "config.vh"

module i_cache (
    input clk,
    input rst,

    
    );
    
endmodule